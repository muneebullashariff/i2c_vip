// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : slave_agt_top.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: slave_agt_top
// Description of the class :
// This class acts like a container to slave agents 
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the slave_agt_top class object
//
// Parameters:
//  name   - instance name of the slave_agt_top
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Function: build_phase
// Creates the slave_agent components 
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------



