module top;

import uvm_pkg::*;
import i2c_pkg::*;

 initial
   begin
     run_test("i2c_test");
   end
endmodule
