// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : master_agt_sequence.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: master_agt_sequence
// Description of the class :
// This class is responsible for generating different stimulus for master
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_agt_sequence class object
//
// Parameters:
//  name   - instance name of the master_agt_sequence
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Task: body
// master_xtn is randomized to get differnet test stimulus
//-----------------------------------------------------------------------------


