// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : i2c_test.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: i2c_test
// Description of the class :
// This class acts like a individual block intended to test the design
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the i2c_test class object
//
// Parameters:
//  name   - instance name of the i2c_test
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: build_phase
// Creates component for environment 
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Task: run_phase
// Starts virtual_sequence on to virtual_sequencer in environment
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------



