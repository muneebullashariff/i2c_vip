// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : scoreboard.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: scoreboard
// Description of the class :
// This class acts like a place to validate data integrity  
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the scoreboard class object
//
// Parameters:
//  name   - instance name of the scoreboard
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: build_phase
// Get the configuration object
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------







