//  ############################################################################
//
//  Licensed to the Apache Software Foundation (ASF) under one
//  or more contributor license agreements.  See the NOTICE file
//  distributed with this work for additional information
//  regarding copyright ownership.  The ASF licenses this file
//  to you under the Apache License, Version 2.0 (the
//  "License"); you may not use this file except in compliance
//  with the License.  You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing,
//  software distributed under the License is distributed on an
//  "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
//  KIND, either express or implied.  See the License for the
//  specific language governing permissions and limitations
//  under the License. 
//
//  ###########################################################################



//-----------------------------------------------------------------------------
// Class: Master_driver
// Description of the class :
// This class drives data to the interface 
//-----------------------------------------------------------------------------

`ifndef master_driver
`define master_driver

class master_driver extends uvm_driver#(master_xtn);
`uvm_component_utils(master_driver)

virtual i2c_intf vif;
master_agent_config mcfg;

//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------

extern function new(string name="master_driver",uvm_component parent);
extern function void build_phase(uvm_phase phase);
extern function void connect_phase(uvm_phase phase);
extern task send_start_bit(master_xtn xtn);
extern task send_slave_address(master_xtn xtn);
extern task send_write_data(master_xtn xtn);
extern task send_stop_bit(master_xtn xtn);
extern task run_phase(uvm_phase phase);

endclass


//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_driver class object
//
// Parameters:
//  name   - instance name of the master_driver
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------


function master_driver::new(string name="master_driver",uvm_component parent);
	super.new(name,parent);
endfunction


//-----------------------------------------------------------------------------
// Function: build_phase
// Creates the required ports
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------


function void master_driver::build_phase(uvm_phase phase);
  if(!uvm_config_db#(master_agent_config)::get(this,"","MASTER_AGENT_CONFIG",mcfg))
   `uvm_fatal("master_driver","COULDNT GET")
endfunction



//-----------------------------------------------------------------------------
// Function: connect_phase
// Connects the master_driver to the required interface
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------


function void master_driver::connect_phase(uvm_phase phase);
vif=mcfg.vif;
endfunction



//-----------------------------------------------------------------------------
// Task: run_phase
// Initiates the main Driving task 
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------

task master_driver::run_phase(uvm_phase phase);

  fork 
    forever
       #(mcfg.clk_period) vif.clk_int=!vif.clk_int;
  join_none

  forever
    begin

 	seq_item_port.get_next_item(req);

	    send_start_bit(req);
	    send_slave_address(req);
	    send_write_data(req);
	    send_stop_bit(req);

	seq_item_port.item_done;

    end
endtask


task master_driver::send_start_bit(master_xtn xtn);
           @(vif.m_drv_cb_ctrl);
	    vif.m_drv_cb_ctrl.sda_int<=xtn.start_bit;
endtask


task master_driver::send_slave_address(master_xtn xtn);
	foreach(xtn.slave_address[i])
	  begin
	    @(vif.m_drv_cb_data);
	    vif.m_drv_cb_data.sda_int<=xtn.slave_address[6-i];
	  end
	    #(mcfg.clk_period/2);
	    vif.sda_int<=1'b1;     //RELEASE SDA LINE SO THAT SLAVE CAN SEND ACK/NACK
endtask


task master_driver::send_write_data(master_xtn xtn);
        foreach(xtn.write_data[i])
	  begin
	    @(vif.m_drv_cb_data);
	     vif.m_drv_cb_data.sda_int<=xtn.write_data[7-i];
	  end
	    #(mcfg.clk_period/2);
	    vif.sda_int<=1'b1;     //RELEASE SDA LINE SO THAT SLAVE CAN SEND ACK/NACK

endtask

task master_driver::send_stop_bit(master_xtn xtn);
           @(vif.m_drv_cb_ctrl);
	    vif.m_drv_cb_ctrl.sda_int<=xtn.stop_bit;
endtask


`endif
