// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : master_agent.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: master_agent
// Description of the class :
// This class acts like a container. 
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_agent class object
//
// Parameters:
//  name   - instance name of the master_agent
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: build_phase
// Creates the components according to is_active value 
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: connect_phase
// Connects master_driver to master_sequencer using TLM Ports if
// is_active==UVM_ACTIVE
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------






