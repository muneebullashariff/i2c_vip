// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : virtual_sequencer.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: virtual_sequencer
// Description of the class :
// This class acts like a container to sequencers of
// master agents and slave agents 
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the virtual_sequencer class object
//
// Parameters:
//  name   - instance name of the virtual_sequencer
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------



