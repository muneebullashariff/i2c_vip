module top;

  initial begin
    $display("Merging concept");
  end
endmodule
