module top;

  initial begin
   $display("VALUE");
  end
endmodule
