// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : slave_agt_sequence.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: slave_agt_sequence
// Description of the class :
// This class is responsible for generating different stimulus for master
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the slave_agt_sequence class object
//
// Parameters:
//  name   - instance name of the slave_agt_sequence
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Task: body
// slave_xtn is randomized to get differnet test stimulus
//-----------------------------------------------------------------------------


