// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : slave_xtn.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: slave_xtn
// Description of the class :
// This class contains variables that would ultimately be provided to
// interface
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the slave_xtn class object
//
// Parameters:
//  name   - instance name of the slave_xtn
//-----------------------------------------------------------------------------


