// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : Master_sequencer.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: Master_sequencer
// Description of the class :
// This class controls the flow of sequence_items between
// master_sequence and master_driver
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_sequencer class object
//
// Parameters:
//  name   - instance name of the master_sequencer
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------

