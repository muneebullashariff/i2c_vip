// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : slave_sequencer.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: slave_sequencer
// Description of the class :
// This class controls the flow of sequence_items between
// slave_sequence and slave_driver
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the slave_sequencer class object
//
// Parameters:
//  name   - instance name of the slave_sequencer
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------

