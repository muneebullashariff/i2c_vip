// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : master_agt_top.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: master_agt_top
// Description of the class :
// This class acts like a container to master agents 
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_agt_top class object
//
// Parameters:
//  name   - instance name of the master_agt_top
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Function: build_phase
// Creates the master_agent components 
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------




