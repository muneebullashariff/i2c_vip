// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : virtual_sequence.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: virtual_sequence
// Description of the class :
// This class is responsible for starting various sequences
// on to respective sequencers 
//-----------------------------------------------------------------------------





//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------



//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the virtual_sequence class object
//
// Parameters:
//  name   - instance name of the virtual_sequence
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Task: body
// master_agt_sequence and slave_agent_sequence is started on 
// respective  sequencers
//-----------------------------------------------------------------------------


