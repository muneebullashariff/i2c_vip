module top;

  initial begin
   $display("VALUE");
   $display("Merging concept");
  end
endmodule
