// ############################################################################
//
// Project : Verification of I2C VIP
//
// File_name : Master_monitor.sv
//
// https://github.com/muneebullashariff/i2c_vip
//
// ############################################################################

//-----------------------------------------------------------------------------
// Class: Master_monitor
// Description of the class :
// This class samples the DUT signals through virtual interface
//-----------------------------------------------------------------------------




//---------------------------------------------
// Externally defined tasks and functions
//---------------------------------------------




//-----------------------------------------------------------------------------
// Constructor: new
// Initializes the master_monitor class object
//
// Parameters:
//  name   - instance name of the master_monitor
//  parent - parent under which this component is created
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: build_phase
// Gets the configuration object
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------






//-----------------------------------------------------------------------------
// Function: connect_phase
// Connects the virtual interface to the interface handle of the monitor
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------





//-----------------------------------------------------------------------------
// Task: run_phase
// Collects the data
//
// Parameters:
//  phase - stores the current phase 
//-----------------------------------------------------------------------------

